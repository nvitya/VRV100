
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity VRV1_365_test_top is
port
(
	FLED 			: out std_logic;
	FKEY 			: in  std_logic;

	BLED 			: out unsigned(4 downto 0);
	BKEY 			: in  unsigned(4 downto 0);

	D7S_SEGMENT : out unsigned(7 downto 0);
   D7S_SEL 		: out unsigned(2 downto 0);

	UART0_TXD_O : out std_logic;
	UART0_RXD_I : in  std_logic := '0';

	SPIM1_SS    : out std_logic;
	SPIM1_SCLK  : out std_logic;
	SPIM1_MOSI  : out std_logic;
	SPIM1_MISO  : in  std_logic;

	JTAG_TCK		: in std_logic;
	JTAG_TDI		: in std_logic;
	JTAG_TDO		: out std_logic;
	JTAG_TMS		: in std_logic;

	DDR3_addr 		: out STD_LOGIC_VECTOR ( 13 downto 0 );
	DDR3_ba 			: out STD_LOGIC_VECTOR ( 2 downto 0 );
	DDR3_cas_n 		: out STD_LOGIC;
	DDR3_ck_n 		: out STD_LOGIC_VECTOR ( 0 to 0 );
	DDR3_ck_p 		: out STD_LOGIC_VECTOR ( 0 to 0 );
	DDR3_cke 		: out STD_LOGIC_VECTOR ( 0 to 0 );
	DDR3_dm 			: out STD_LOGIC_VECTOR ( 1 downto 0 );
	DDR3_dq 			: inout STD_LOGIC_VECTOR ( 15 downto 0 );
	DDR3_dqs_n 		: inout STD_LOGIC_VECTOR ( 1 downto 0 );
	DDR3_dqs_p 		: inout STD_LOGIC_VECTOR ( 1 downto 0 );
	DDR3_odt 		: out STD_LOGIC_VECTOR ( 0 to 0 );
	DDR3_ras_n 		: out STD_LOGIC;
	DDR3_reset_n 	: out STD_LOGIC;
	DDR3_we_n 		: out STD_LOGIC;

	CLKIN_50 	: in std_logic -- 50 MHz clock
);
end entity;

architecture behavioral of VRV1_365_test_top
is
	signal CLKCNT : unsigned(31 downto 0);
	signal CLK : std_logic;

	signal RESET 		: std_logic;
	signal RESET_N    : std_ulogic;

	signal CLK_100_PLL	: std_logic;
	signal CLK_100_AXI	: std_logic;  -- generated by the DDR3 controller

	signal GPIO_OUT 		: std_logic_vector(31 downto 0);

	signal GPIOA_IO      : std_logic_vector(31 downto 0);
	signal GPIOB_IO      : std_logic_vector(31 downto 0);

	signal AXI_AW_VALID 				: std_logic;
	signal AXI_AW_READY 				: std_logic;
	signal AXI_AW_PAYLOAD_ADDR 	: std_logic_vector(27 downto 0);
	signal AXI_AW_PAYLOAD_ID 		: std_logic_vector( 3 downto 0);
	signal AXI_AW_PAYLOAD_LEN 		: std_logic_vector( 7 downto 0);
	signal AXI_AW_PAYLOAD_SIZE 	: std_logic_vector( 2 downto 0);
	signal AXI_AW_PAYLOAD_BURST 	: std_logic_vector( 1 downto 0);
	signal AXI_AW_PAYLOAD_LOCK 	: std_logic_vector( 0 downto 0);
	signal AXI_AW_PAYLOAD_CACHE 	: std_logic_vector( 3 downto 0);
	signal AXI_AW_PAYLOAD_QOS 		: std_logic_vector( 3 downto 0);
	signal AXI_AW_PAYLOAD_PROT 	: std_logic_vector( 2 downto 0);
	signal AXI_W_VALID 				: std_logic;
	signal AXI_W_READY 				: std_logic;
	signal AXI_W_PAYLOAD_DATA 		: std_logic_vector(31 downto 0);
	signal AXI_W_PAYLOAD_STRB 		: std_logic_vector( 3 downto 0);
	signal AXI_W_PAYLOAD_LAST 		: std_logic;
	signal AXI_B_VALID 				: std_logic;
	signal AXI_B_READY 				: std_logic;
	signal AXI_B_PAYLOAD_ID 		: std_logic_vector( 3 downto 0);
	signal AXI_B_PAYLOAD_RESP 		: std_logic_vector( 1 downto 0);
	signal AXI_AR_VALID 				: std_logic;
	signal AXI_AR_READY 				: std_logic;
	signal AXI_AR_PAYLOAD_ADDR 	: std_logic_vector(27 downto 0);
	signal AXI_AR_PAYLOAD_ID 		: std_logic_vector( 3 downto 0);
	signal AXI_AR_PAYLOAD_LEN 		: std_logic_vector( 7 downto 0);
	signal AXI_AR_PAYLOAD_SIZE 	: std_logic_vector( 2 downto 0);
	signal AXI_AR_PAYLOAD_BURST 	: std_logic_vector( 1 downto 0);
	signal AXI_AR_PAYLOAD_LOCK 	: std_logic_vector( 0 downto 0);
	signal AXI_AR_PAYLOAD_CACHE 	: std_logic_vector( 3 downto 0);
	signal AXI_AR_PAYLOAD_QOS 		: std_logic_vector( 3 downto 0);
	signal AXI_AR_PAYLOAD_PROT 	: std_logic_vector( 2 downto 0);
	signal AXI_R_VALID 				: std_logic;
	signal AXI_R_READY 				: std_logic;
	signal AXI_R_PAYLOAD_DATA 		: std_logic_vector(31 downto 0);
	signal AXI_R_PAYLOAD_ID 		: std_logic_vector( 3 downto 0);
	signal AXI_R_PAYLOAD_RESP 		: std_logic_vector( 1 downto 0);
	signal AXI_R_PAYLOAD_LAST 		: std_logic;

	signal APB_PADDR		: std_logic_vector(19 downto 0);
	signal APB_PSEL		: std_logic;
	signal APB_PENABLE	: std_logic;
	signal APB_PREADY		: std_logic;
	signal APB_PWRITE		: std_logic;
	signal APB_PWDATA		: std_logic_vector(31 downto 0);
	signal APB_PRDATA		: std_logic_vector(31 downto 0);
	signal APB_PSLVERROR	: std_logic;

   component clock_pll
   port
   (
     clk_out1  : out    std_logic;
     clk_in1   : in     std_logic
   );
   end component;

begin
	RESET_N <= FKEY;
	RESET <= not RESET_N;

	CLK 	 <= CLK_100_AXI;

	FLED <= GPIOA_IO(0);

   clockgen : component clock_pll
   port map
   (
      clk_out1 => CLK_100_PLL,
      clk_in1  => CLKIN_50
   );

   ext_ram : entity work.ddr3_ram
   port map
   (
		AXI_awvalid 	=> AXI_AW_VALID,
		AXI_awready 	=> AXI_AW_READY,
		AXI_awaddr 		=> AXI_AW_PAYLOAD_ADDR,
		AXI_awid 		=> AXI_AW_PAYLOAD_ID,
		AXI_awlen 		=> AXI_AW_PAYLOAD_LEN,
		AXI_awsize 		=>	AXI_AW_PAYLOAD_SIZE,
		AXI_awburst 	=> AXI_AW_PAYLOAD_BURST,
		AXI_awlock 		=> AXI_AW_PAYLOAD_LOCK(0),
		AXI_awcache 	=> AXI_AW_PAYLOAD_CACHE,
		AXI_awqos 		=> AXI_AW_PAYLOAD_QOS,
		AXI_awprot 		=> AXI_AW_PAYLOAD_PROT,
		AXI_wvalid 		=> AXI_W_VALID,
		AXI_wready 		=> AXI_W_READY,
		AXI_wdata 		=> AXI_W_PAYLOAD_DATA,
		AXI_wstrb 		=> AXI_W_PAYLOAD_STRB,
		AXI_wlast 		=> AXI_W_PAYLOAD_LAST,
		AXI_bvalid 		=> AXI_B_VALID,
		AXI_bready 		=> AXI_B_READY,
		AXI_bid 			=> AXI_B_PAYLOAD_ID,
		AXI_bresp 		=> AXI_B_PAYLOAD_RESP,
		AXI_arvalid		=> AXI_AR_VALID,
		AXI_arready 	=> AXI_AR_READY,
		AXI_araddr 		=> AXI_AR_PAYLOAD_ADDR,
		AXI_arid 		=> AXI_AR_PAYLOAD_ID,
		AXI_arlen 		=> AXI_AR_PAYLOAD_LEN,
		AXI_arsize 		=> AXI_AR_PAYLOAD_SIZE,
		AXI_arburst 	=> AXI_AR_PAYLOAD_BURST,
		AXI_arlock 		=> AXI_AR_PAYLOAD_LOCK(0),
		AXI_arcache 	=> AXI_AR_PAYLOAD_CACHE,
		AXI_arqos 		=> AXI_AR_PAYLOAD_QOS,
		AXI_arprot 		=> AXI_AR_PAYLOAD_PROT,
		AXI_rvalid 		=> AXI_R_VALID,
		AXI_rready 		=> AXI_R_READY,
		AXI_rdata 		=> AXI_R_PAYLOAD_DATA,
		AXI_rid 			=> AXI_R_PAYLOAD_ID,
		AXI_rresp 		=> AXI_R_PAYLOAD_RESP,
		AXI_rlast 		=> AXI_R_PAYLOAD_LAST,

		DDR3_addr 		=> DDR3_addr,
		DDR3_ba 			=> DDR3_ba,
		DDR3_cas_n 		=> DDR3_cas_n,
		DDR3_ck_n 		=> DDR3_ck_n,
		DDR3_ck_p 		=> DDR3_ck_p,
		DDR3_cke 		=> DDR3_cke,
		DDR3_dm 			=> DDR3_dm,
		DDR3_dq 			=> DDR3_dq,
		DDR3_dqs_n 		=> DDR3_dqs_n,
		DDR3_dqs_p 		=> DDR3_dqs_p,
		DDR3_odt 		=> DDR3_odt,
		DDR3_ras_n 		=> DDR3_ras_n,
		DDR3_reset_n 	=> DDR3_reset_n,
		DDR3_we_n 		=> DDR3_we_n,

		AXI_CLK_OUT 	=> CLK_100_AXI,
		CLK_100_IN 		=> CLK_100_PLL,
		RESET_N 			=> RESET_N
   );

	u0 : entity work.VRV1_365_vhdl
	port map
	(
		GPIOA_IO					=>	GPIOA_IO,
		GPIOB_IO					=>	GPIOB_IO,

		UART1_TXD_O 			=> UART0_TXD_O,
		UART1_RXD_I 			=> UART0_RXD_I,

		UART2_TXD_O 			=> open,
		UART2_RXD_I 			=> '1',

		SPIM1_SS(0)   			=> SPIM1_SS,
		SPIM1_SS(3 downto 1) => open,
		SPIM1_SCLK  			=> SPIM1_SCLK,
		SPIM1_MOSI  			=> SPIM1_MOSI,
		SPIM1_MISO  			=> SPIM1_MISO,

		SPIM2_SS    			=> open,
		SPIM2_SCLK  			=> open,
		SPIM2_MOSI  			=> open,
		SPIM2_MISO  			=> '0',

		AXI_AW_VALID 				=> AXI_AW_VALID,
		AXI_AW_READY 				=> AXI_AW_READY,
		AXI_AW_PAYLOAD_ADDR 	   => AXI_AW_PAYLOAD_ADDR,
		AXI_AW_PAYLOAD_ID 		=> AXI_AW_PAYLOAD_ID,
		AXI_AW_PAYLOAD_LEN 		=> AXI_AW_PAYLOAD_LEN,
		AXI_AW_PAYLOAD_SIZE 	   => AXI_AW_PAYLOAD_SIZE,
		AXI_AW_PAYLOAD_BURST 	=> AXI_AW_PAYLOAD_BURST,
		AXI_AW_PAYLOAD_LOCK 	   => AXI_AW_PAYLOAD_LOCK,
		AXI_AW_PAYLOAD_CACHE 	=> AXI_AW_PAYLOAD_CACHE,
		AXI_AW_PAYLOAD_QOS 		=> AXI_AW_PAYLOAD_QOS,
		AXI_AW_PAYLOAD_PROT 		=> AXI_AW_PAYLOAD_PROT,
		AXI_W_VALID 				=> AXI_W_VALID,
		AXI_W_READY 				=> AXI_W_READY,
		AXI_W_PAYLOAD_DATA 		=> AXI_W_PAYLOAD_DATA,
		AXI_W_PAYLOAD_STRB 		=> AXI_W_PAYLOAD_STRB,
		AXI_W_PAYLOAD_LAST 		=> AXI_W_PAYLOAD_LAST,
		AXI_B_VALID 				=> AXI_B_VALID,
		AXI_B_READY 				=> AXI_B_READY,
		AXI_B_PAYLOAD_ID 			=> AXI_B_PAYLOAD_ID,
		AXI_B_PAYLOAD_RESP 		=> AXI_B_PAYLOAD_RESP,
		AXI_AR_VALID 				=> AXI_AR_VALID,
		AXI_AR_READY 				=> AXI_AR_READY,
		AXI_AR_PAYLOAD_ADDR 		=> AXI_AR_PAYLOAD_ADDR,
		AXI_AR_PAYLOAD_ID 		=> AXI_AR_PAYLOAD_ID,
		AXI_AR_PAYLOAD_LEN 		=> AXI_AR_PAYLOAD_LEN,
		AXI_AR_PAYLOAD_SIZE 		=> AXI_AR_PAYLOAD_SIZE,
		AXI_AR_PAYLOAD_BURST 	=> AXI_AR_PAYLOAD_BURST,
		AXI_AR_PAYLOAD_LOCK 		=> AXI_AR_PAYLOAD_LOCK,
		AXI_AR_PAYLOAD_CACHE 	=> AXI_AR_PAYLOAD_CACHE,
		AXI_AR_PAYLOAD_QOS 		=> AXI_AR_PAYLOAD_QOS,
		AXI_AR_PAYLOAD_PROT 		=> AXI_AR_PAYLOAD_PROT,
		AXI_R_VALID 				=> AXI_R_VALID,
		AXI_R_READY 				=> AXI_R_READY,
		AXI_R_PAYLOAD_DATA 		=> AXI_R_PAYLOAD_DATA,
		AXI_R_PAYLOAD_ID 			=> AXI_R_PAYLOAD_ID,
		AXI_R_PAYLOAD_RESP 		=> AXI_R_PAYLOAD_RESP,
		AXI_R_PAYLOAD_LAST 		=> AXI_R_PAYLOAD_LAST,

		JTAG_TMS            	=> JTAG_TMS,
		JTAG_TDI            	=> JTAG_TDI,
		JTAG_TDO            	=> JTAG_TDO,
		JTAG_TCK            	=> JTAG_TCK,

		APB_PADDR				=> APB_PADDR,
		APB_PSEL					=> APB_PSEL,
		APB_PENABLE				=> APB_PENABLE,
		APB_PREADY				=> APB_PREADY,
		APB_PWRITE				=> APB_PWRITE,
		APB_PWDATA				=> APB_PWDATA,
		APB_PRDATA				=> APB_PRDATA,
		APB_PSLVERROR			=> APB_PSLVERROR,

		CLK_100	            => CLK,
		RESET						=> RESET
	);

	periph : entity work.apb_periph
	port map
	(
		APB_PADDR		=> APB_PADDR,
		APB_PSEL			=> APB_PSEL,
		APB_PENABLE		=> APB_PENABLE,
		APB_PREADY		=> APB_PREADY,
		APB_PWRITE		=> APB_PWRITE,
		APB_PWDATA		=> APB_PWDATA,
		APB_PRDATA		=> APB_PRDATA,
		APB_PSLVERROR	=> APB_PSLVERROR,

		GPIO_OUT			=> GPIO_OUT,
		GPIO_IN			=> std_logic_vector(CLKCNT(31 downto 0)),

		RESET     		=> RESET,
		CLK		 		=> CLK
	);

	process (CLK)
	begin
	 if rising_edge(CLK)
	 then
		CLKCNT <= CLKCNT + 1;
	 end if;
	end process;

end architecture;
